-- -------------------------------------------------------------------------------------------------
-- Copyright (c) Lukas Vik. All rights reserved.
-- Copyright (c) DESY
--
-- Original file is part of the tsfpga project.
-- https://tsfpga.com
-- https://gitlab.com/tsfpga/tsfpga
--
-- Modified file is part of the hdl_modules fork
-- https://github.com/nicdes/hdl-modules
-- Changes:
-- * added async reset logic
-- * added axi write strobe handling (big or little endian)
-- * refactoring with double buffer for atomic read/write.
-- * regs_up_valid
-- -------------------------------------------------------------------------------------------------
-- General register file controlled over AXI-Lite.
--
-- Will respond with ``SLVERR`` on the ``R`` channel when attempting to read a register that
--
-- 1. Does not exists (``ARADDR`` out of range), or
-- 2. Is not of a register type that can be read by the bus (e.g. write only).
--
-- Similarly it will respond with ``SLVERR`` on the ``B`` channel attempting to write a
-- register that
--
-- 1. Does not exists (``AWADDR`` out of range), or
-- 2. Is not of a register type that can be written by the bus (e.g. read only).
--
-- Both cases are handled cleanly without stalling or hanging the AXI-Lite bus.
--
-- The ``regs`` and ``default_values`` generics are designed to get their values
-- from a package generated by the ``hdl_registers`` VHDL generator:
-- :py:class:`RegisterVhdlGenerator <hdl_registers.register_vhdl_generator.RegisterVhdlGenerator>`.
-- The values can be constructed by hand as well, of course.
-- -------------------------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library common;
use common.addr_pkg.all;

library axi;
use axi.axi_pkg.all;
use axi.axi_lite_pkg.all;

use work.reg_file_pkg.all;

entity axi_lite_reg_file is
  generic (
    regs           : reg_definition_vec_t;
    default_values : reg_vec_t(regs'range) := (others => (others => '0'));
    use_wstrb      : boolean               := false;
    -- If 'big' wstrb(0) qualifies the most significant byte.  If 'small', the
    -- least significant.
    big_endian     : boolean               := true  -- true for big, false for little
    );
  port (
    rst_n            : in  std_ulogic;
    clk              : in  std_logic;
    --# {{}}
    --# Register control bus
    axi_lite_m2s     : in  axi_lite_m2s_t;
    axi_lite_s2m     : out axi_lite_s2m_t;
    --# {{}}
    -- Register values
    -- Assert regs_up_slverr to force a slave error AXI read response.
    -- A slave error AXI response is sent anyway if reading from a unknown
    -- address.
    regs_down        : out reg_vec_t(regs'range);
    regs_up          : in  reg_vec_t(regs'range)         := default_values;
    regs_up_valid    : in  std_ulogic_vector(regs'range) := (others => '1');
    regs_up_ready    : out std_ulogic_vector(regs'range) := (others => '0');
    regs_up_slverr   : in  std_ulogic_vector(regs'range) := (others => '0');
    regs_down_slverr : in  std_ulogic_vector(regs'range) := (others => '0');
    --# {{}}
    -- Each bit is pulsed for one cycle when the corresponding register is read/written.
    -- For read, the bit is asserted the exact same cycle as the AXI-Lite R transaction occurs.
    -- For write, the bit is asserted the cycle after the AXI-Lite W transaction occurs, so that
    -- 'regs_down' is updated with the new value.
    reg_was_read     : out std_logic_vector(regs'range);
    reg_was_written  : out std_logic_vector(regs'range);
    reg_down_strb    : out std_ulogic_vector(axi_lite_w_strb_sz-1 downto 0)
    );
end entity;

architecture a of axi_lite_reg_file is

  constant addr_and_mask_vec : addr_and_mask_vec_t := to_addr_and_mask_vec(regs);

  constant invalid_addr : integer := regs'length;
  subtype decoded_idx_t is integer range 0 to invalid_addr;

  signal s_reg_values_read_buf  : reg_vec_t(regs'range);
  signal s_reg_values_write_buf : reg_vec_t(regs'range);

  signal s_reg_being_read              : std_ulogic_vector(regs'range);
  signal s_reg_was_written             : std_ulogic_vector(regs'range);
  signal s_atomic_read, s_atomic_write : std_ulogic_vector(regs'range);

  function is_atomic (
    constant idx : integer range regs'range)
    return boolean is
  begin
    for i in regs'range loop
      if i <= idx then
        if regs(i).atomic_lock /= 0 then
          if idx <= i + regs(i).atomic_lock then
            return true;
          end if;
        end if;
      end if;
    end loop;

    return false;
  end function is_atomic;

begin

  -- s_atomic_read and s_atomic_write from
  -- s_reg_begin_read and s_reg_was_written
  -- Note: this is fine for synthesis because atomic_lock indexes are
  -- static.
  atomic_double_buffer_block : block is
  begin
    atomic_read_proc : process (all) is
    begin
      s_atomic_read <= (others => '0');
      for idx in regs'range loop
        if s_reg_being_read(idx) then
          if is_atomic_segment_start(regs(idx)) then
            s_atomic_read(idx to idx + regs(idx).atomic_lock) <= (others => '1');
          end if;
        end if;
      end loop;
    end process atomic_read_proc;

    atomic_write_proc : process (all) is
    begin
      s_atomic_write <= (others => '0');

      for idx in regs'range loop
        if s_reg_was_written(idx) then
          if is_atomic_segment_end(regs(idx)) then
            s_atomic_write(idx + regs(idx).atomic_lock to idx) <= (others => '1');
          end if;
        end if;
      end loop;
    end process atomic_write_proc;
  end block atomic_double_buffer_block;

  read_block : block
    type read_state_t is (ar, atomic_read, r);
    signal read_state : read_state_t;
  begin

    read_process : process (clk, rst_n) is
      variable v_data        : reg_t;
      variable v_read_idx    : integer range regs'range;
      variable v_decoded_idx : decoded_idx_t;

      -- An address transaction has occured and the address points to a valid
      -- read register
      function is_valid_read_address (
        idx : integer) return boolean is
      begin
        return (
          idx /= invalid_addr and
          is_read_type(regs(idx).reg_type));
      end function;

      -- purpose: set axi read data and read response. If address is valid
      -- response is okay, else slverr.
      procedure set_axi_response (
        idx  : natural;
        data : reg_t
        ) is
      begin
        if is_valid_read_address(idx) and regs_up_slverr(idx) = '0' then
          axi_lite_s2m.read.r.resp <= axi_resp_okay;
          axi_lite_s2m.read.r.data <= data;
        else
          axi_lite_s2m.read.r.resp <= axi_resp_slverr;
          axi_lite_s2m.read.r.data <= (others => '-');
        end if;
      end procedure set_axi_response;

    begin
      if not rst_n then
        axi_lite_s2m.read <= (
          ar => (ready => '1'),
          r  => axi_lite_s2m_r_init);
        reg_was_read     <= (others => '0');
        regs_up_ready    <= (others => '0');
        s_reg_being_read <= (others => '0');

        read_state    <= ar;
        v_data        := (others => '-');
        v_decoded_idx := invalid_addr;
        v_read_idx    := 0;

        s_reg_values_read_buf <= (others => (others => '-'));
        for idx in regs'range loop
          if is_fabric_gives_value_type(regs(idx).reg_type) and is_atomic(idx) then
            s_reg_values_read_buf(idx) <= (others => '0');
          end if;
        end loop;
      elsif rising_edge(clk) then

        axi_lite_s2m.read <= axi_lite_read_s2m_init;

        reg_was_read <= (others => '0');
        v_data       := (others => '-');

        case read_state is
          when ar =>
            v_read_idx    := 0;
            v_decoded_idx := invalid_addr;

            axi_lite_s2m.read.ar.ready <= '1';
            regs_up_ready              <= (others => '0');
            s_reg_being_read           <= (others => '-');

            if axi_lite_m2s.read.ar.valid and axi_lite_s2m.read.ar.ready then
              axi_lite_s2m.read.ar.ready <= '0';
              v_decoded_idx              := decode(axi_lite_m2s.read.ar.addr, addr_and_mask_vec);
              if v_decoded_idx /= invalid_addr then
                v_read_idx := v_decoded_idx;
              end if;
              s_reg_being_read(v_read_idx) <= '1';

              if is_atomic(v_read_idx) then
                read_state <= atomic_read;
              else
                read_state <= r;
              end if;
            end if;

          when atomic_read =>
            -- Transfer data to to the double buffer from regs_up if fabric
            -- gives value.  This is done here to easy timing on the decoder
            -- state (ar).
            read_state <= r;

            for idx in regs'range loop
              if s_atomic_read(idx) then
                if is_fabric_gives_value_type(regs(idx).reg_type) then
                  if regs_up_valid(idx) then
                    s_reg_values_read_buf(idx) <= regs_up(idx);
                  else
                    read_state <= atomic_read;
                  end if;
                end if;
              end if;
            end loop;

          when r =>

            axi_lite_s2m.read.r.valid <= '1';
            regs_up_ready(v_read_idx) <= '1';

            if is_fabric_gives_value_type(regs(v_read_idx).reg_type) then
              if is_atomic(v_read_idx) then
                v_data := s_reg_values_read_buf(v_read_idx);
              else
                if not regs_up_valid(v_read_idx) then
                  -- hold off transaction if regs_up_valid(idx) is
                  -- deasserted.  This is done for atomic registers in
                  -- the atomic_read state.
                  axi_lite_s2m.read.r.valid <= '0';
                else
                  v_data := regs_up(v_read_idx);
                end if;
              end if;
            else
              v_data := regs_down(v_read_idx);
            end if;

            set_axi_response(v_read_idx, v_data);

            if axi_lite_m2s.read.r.ready and axi_lite_s2m.read.r.valid then
              axi_lite_s2m.read.r.valid  <= '0';
              axi_lite_s2m.read.ar.ready <= '1';
              regs_up_ready              <= (others => '0');

              if is_valid_read_address(v_read_idx) then
                if is_atomic(v_read_idx) then
                  if is_atomic_segment_end(regs(v_read_idx)) then
                    reg_was_read(v_read_idx) <= '1';
                  end if;
                else
                  reg_was_read(v_read_idx) <= '1';
                end if;
              end if;

              read_state <= ar;
            end if;

        end case;

      end if;
    end process;
  end block;

  write_block : block
    type write_state_t is (aw, w, atomic_write, b);
    signal write_state : write_state_t;
  begin

    write_process : process (clk, rst_n) is
      variable v_byte_idx    : integer range 0 to axi_lite_w_strb_sz-1;
      variable v_decoded_idx : decoded_idx_t;
      variable v_write_idx   : integer range regs'range;
      variable v_data        : reg_t;

      -- An address transaction has occured and the address points to a valid
      -- write register
      function is_valid_write_address (
        idx : integer) return boolean is
      begin
        return idx /= invalid_addr and
          is_write_type(regs(idx).reg_type);
      end function;

      -- purpose: set axi write response. If address is valid response is okay,
      -- else slverr.
      procedure set_axi_response (
        idx : natural
        ) is
      begin
        axi_lite_s2m.write.b.valid <= '1';
        if is_valid_write_address(idx) and regs_down_slverr(idx) = '0' then
          axi_lite_s2m.write.b.resp <= axi_resp_okay;
        else
          axi_lite_s2m.write.b.resp <= axi_resp_slverr;
        end if;
      end procedure set_axi_response;

    begin
      if not rst_n then
        axi_lite_s2m.write <= axi_lite_write_s2m_init;
        reg_was_written    <= (others => '0');
        s_reg_was_written  <= (others => '0');
        write_state        <= aw;
        v_decoded_idx      := invalid_addr;
        v_write_idx        := 0;
        v_data             := (others => '-');

        regs_down     <= default_values;
        reg_down_strb <= (others => '0');

        s_reg_values_write_buf <= (others => (others => '-'));
        for idx in regs'range loop
          if is_write_type(regs(idx).reg_type) then
            if is_atomic(idx) then
              s_reg_values_write_buf(idx) <= (others => '0');
            end if;
          end if;
        end loop;
      elsif rising_edge(clk) then

        axi_lite_s2m.write <= axi_lite_write_s2m_init;
        reg_down_strb      <= (others => '0');
        reg_was_written    <= (others => '0');
        s_reg_was_written  <= (others => '0');
        v_data             := (others => '-');

        -- clear write pulse registers
        for idx in regs'range loop
          if is_write_pulse_type(regs(idx).reg_type) then
            regs_down(idx) <= (others => '0');
          end if;
        end loop;

        case write_state is
          when aw =>
            v_write_idx   := 0;
            v_decoded_idx := invalid_addr;

            axi_lite_s2m.write.aw.ready <= '1';
            if axi_lite_m2s.write.aw.valid and axi_lite_s2m.write.aw.ready then
              axi_lite_s2m.write.aw.ready <= '0';

              v_decoded_idx := decode(axi_lite_m2s.write.aw.addr, addr_and_mask_vec);
              if v_decoded_idx /= invalid_addr then
                v_write_idx := v_decoded_idx;
              end if;
              axi_lite_s2m.write.w.ready <= '1';
              write_state                <= w;
            end if;

          when w =>
            axi_lite_s2m.write.w.ready <= '1';
            if axi_lite_m2s.write.w.valid and axi_lite_s2m.write.w.ready then
              axi_lite_s2m.write.w.ready <= '0';

              if is_valid_write_address(v_write_idx) then
                s_reg_was_written(v_write_idx) <= '1';

                if use_wstrb then
                  if is_atomic(v_write_idx) then
                    v_data := s_reg_values_write_buf(v_write_idx);
                  else
                    v_data := regs_down(v_write_idx);
                  end if;

                  for i in axi_lite_m2s.write.w.strb'range loop
                    if axi_lite_m2s.write.w.strb(i) then

                      if not big_endian then
                        v_byte_idx := i;
                      else
                        v_byte_idx := axi_lite_w_strb_sz-i-1;
                      end if;

                      v_data(
                        (v_byte_idx+1)*8-1 downto v_byte_idx*8) := axi_lite_m2s.write.w.data((v_byte_idx+1)*8-1 downto v_byte_idx*8);
                    end if;
                  end loop;

                else
                  -- not using write strobe => write all bytes.
                  v_data := axi_lite_m2s.write.w.data;
                end if;

              end if;

              if is_atomic(v_write_idx) then
                -- write at next state
                write_state                         <= atomic_write;
                s_reg_values_write_buf(v_write_idx) <= v_data;
              else
                write_state <= b;

                regs_down(v_write_idx)       <= v_data;
                reg_was_written(v_write_idx) <= '1';
                reg_down_strb                <= axi_lite_m2s.write.w.strb;
              end if;

            else
              write_state <= b;
            end if;

          when atomic_write =>
            -- Transfer data from s_reg_values_write_buf to regs_down.
            write_state <= b;

            if is_valid_write_address(v_write_idx) then
              if is_atomic(v_write_idx) then
                for idx in regs'range loop
                  if s_atomic_write(idx) then
                    regs_down(idx) <= s_reg_values_write_buf(idx);

                    if is_atomic_segment_end(regs(idx)) then
                      reg_was_written(v_write_idx) <= '1';
                      reg_down_strb                <= axi_lite_m2s.write.w.strb;
                    end if;
                  end if;
                end loop;
              end if;
            end if;

          when b =>
            axi_lite_s2m.write.b.valid <= '1';
            set_axi_response(v_write_idx);
            if axi_lite_m2s.write.b.ready and axi_lite_s2m.write.b.valid then
              axi_lite_s2m.write.aw.ready <= '1';
              axi_lite_s2m.write.b.valid  <= '0';
              write_state                 <= aw;

            end if;
        end case;

      end if;
    end process;
  end block;

end architecture;
